-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"9c080b0b",
    10 => x"0bbda008",
    11 => x"0b0b0bbd",
    12 => x"a4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bda40c0b",
    16 => x"0b0bbda0",
    17 => x"0c0b0b0b",
    18 => x"bd9c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb1cc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bd9c7080",
    57 => x"c7cc278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188c804",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbdac0c",
    65 => x"9f0bbdb0",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bdb008ff",
    69 => x"05bdb00c",
    70 => x"bdb00880",
    71 => x"25eb38bd",
    72 => x"ac08ff05",
    73 => x"bdac0cbd",
    74 => x"ac088025",
    75 => x"d738800b",
    76 => x"bdb00c80",
    77 => x"0bbdac0c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbdac08",
    97 => x"258f3882",
    98 => x"bd2dbdac",
    99 => x"08ff05bd",
   100 => x"ac0c82ff",
   101 => x"04bdac08",
   102 => x"bdb00853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bdac08a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bdb0",
   111 => x"088105bd",
   112 => x"b00cbdb0",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbdb00c",
   116 => x"bdac0881",
   117 => x"05bdac0c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bd",
   122 => x"b0088105",
   123 => x"bdb00cbd",
   124 => x"b008a02e",
   125 => x"0981068e",
   126 => x"38800bbd",
   127 => x"b00cbdac",
   128 => x"088105bd",
   129 => x"ac0c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbdb4",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbdb40c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bd",
   169 => x"b4088407",
   170 => x"bdb40c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb8ac",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bdb40852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bd9c0c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"92710c86",
   219 => x"a42d8271",
   220 => x"0c028405",
   221 => x"0d0402dc",
   222 => x"050d7a54",
   223 => x"800bbdbc",
   224 => x"08f80c89",
   225 => x"1580f52d",
   226 => x"8a1680f5",
   227 => x"2d718280",
   228 => x"29058817",
   229 => x"80f52d70",
   230 => x"84808029",
   231 => x"12f40c52",
   232 => x"555659a4",
   233 => x"0bec0c73",
   234 => x"52bdb851",
   235 => x"a8ea2dbd",
   236 => x"9c08792e",
   237 => x"80eb38bd",
   238 => x"bc0879ff",
   239 => x"12565956",
   240 => x"73792e8b",
   241 => x"38811874",
   242 => x"812a5558",
   243 => x"73f738f7",
   244 => x"18588159",
   245 => x"80762580",
   246 => x"c8387752",
   247 => x"7351848b",
   248 => x"2dbe8452",
   249 => x"bdb851ab",
   250 => x"a92dbd9c",
   251 => x"08802e9a",
   252 => x"38be8457",
   253 => x"83fc5576",
   254 => x"70840558",
   255 => x"08e80cfc",
   256 => x"15557480",
   257 => x"25f13888",
   258 => x"9104bd9c",
   259 => x"08598480",
   260 => x"56bdb851",
   261 => x"aafb2dfc",
   262 => x"80168115",
   263 => x"555687d4",
   264 => x"0486b72d",
   265 => x"840bec0c",
   266 => x"78802e8d",
   267 => x"38b8b051",
   268 => x"91902d8f",
   269 => x"932d88bf",
   270 => x"04baec51",
   271 => x"91902d78",
   272 => x"bd9c0c02",
   273 => x"a4050d04",
   274 => x"02e0050d",
   275 => x"8055840b",
   276 => x"ec0c8ef4",
   277 => x"2d8bde2d",
   278 => x"81f82d9f",
   279 => x"df2dbd9c",
   280 => x"08752e82",
   281 => x"e4388c0b",
   282 => x"ec0cb6ec",
   283 => x"52bdb851",
   284 => x"a8ea2dbd",
   285 => x"9c08752e",
   286 => x"80e538bd",
   287 => x"bc0875ff",
   288 => x"12565956",
   289 => x"73752e8b",
   290 => x"38811874",
   291 => x"812a5558",
   292 => x"73f738f7",
   293 => x"18588076",
   294 => x"2580c438",
   295 => x"77527351",
   296 => x"848b2dbe",
   297 => x"8452bdb8",
   298 => x"51aba92d",
   299 => x"bd9c0880",
   300 => x"2e9a38be",
   301 => x"845783fc",
   302 => x"55767084",
   303 => x"055808e8",
   304 => x"0cfc1555",
   305 => x"748025f1",
   306 => x"3889cf04",
   307 => x"848056bd",
   308 => x"b851aafb",
   309 => x"2dfc8016",
   310 => x"81155556",
   311 => x"899604bd",
   312 => x"bc08f80c",
   313 => x"86b72d84",
   314 => x"0bec0c86",
   315 => x"f651b1c3",
   316 => x"2db8b051",
   317 => x"91902d8f",
   318 => x"932d8bea",
   319 => x"2d91a02d",
   320 => x"b8d00b80",
   321 => x"f52d7082",
   322 => x"2b9c06b8",
   323 => x"c40b80f5",
   324 => x"2d830671",
   325 => x"07b8dc0b",
   326 => x"80f52d70",
   327 => x"852ba006",
   328 => x"b8e80b80",
   329 => x"f52d7086",
   330 => x"2b80c006",
   331 => x"74730707",
   332 => x"b8f40b80",
   333 => x"f52d7087",
   334 => x"2b818006",
   335 => x"b9800b80",
   336 => x"f52d7088",
   337 => x"2b828006",
   338 => x"74730707",
   339 => x"b98c0b80",
   340 => x"f52d7089",
   341 => x"2b848006",
   342 => x"b9980b80",
   343 => x"f52d708a",
   344 => x"2b888006",
   345 => x"74730707",
   346 => x"b9a40b80",
   347 => x"f52d708b",
   348 => x"2b908006",
   349 => x"b9b00b80",
   350 => x"f52d708c",
   351 => x"2ba08006",
   352 => x"74730707",
   353 => x"b9bc0b80",
   354 => x"f52d708d",
   355 => x"2b81c080",
   356 => x"06b9c80b",
   357 => x"80f52d70",
   358 => x"8f2b8280",
   359 => x"80067473",
   360 => x"0707fc0c",
   361 => x"54545454",
   362 => x"54545454",
   363 => x"54545454",
   364 => x"54545454",
   365 => x"5b545257",
   366 => x"54548653",
   367 => x"bd9c0883",
   368 => x"38845372",
   369 => x"ec0c89fa",
   370 => x"04800bbd",
   371 => x"9c0c02a0",
   372 => x"050d0471",
   373 => x"980c04ff",
   374 => x"b008bd9c",
   375 => x"0c04810b",
   376 => x"ffb00c04",
   377 => x"800bffb0",
   378 => x"0c0402f4",
   379 => x"050d8cec",
   380 => x"04bd9c08",
   381 => x"81f02e09",
   382 => x"81068938",
   383 => x"810bbbd0",
   384 => x"0c8cec04",
   385 => x"bd9c0881",
   386 => x"e02e0981",
   387 => x"06893881",
   388 => x"0bbbd40c",
   389 => x"8cec04bd",
   390 => x"9c0852bb",
   391 => x"d408802e",
   392 => x"8838bd9c",
   393 => x"08818005",
   394 => x"5271842c",
   395 => x"728f0653",
   396 => x"53bbd008",
   397 => x"802e9938",
   398 => x"728429bb",
   399 => x"90057213",
   400 => x"81712b70",
   401 => x"09730806",
   402 => x"730c5153",
   403 => x"538ce204",
   404 => x"728429bb",
   405 => x"90057213",
   406 => x"83712b72",
   407 => x"0807720c",
   408 => x"5353800b",
   409 => x"bbd40c80",
   410 => x"0bbbd00c",
   411 => x"bdc4518d",
   412 => x"ed2dbd9c",
   413 => x"08ff24fe",
   414 => x"f838800b",
   415 => x"bd9c0c02",
   416 => x"8c050d04",
   417 => x"02f8050d",
   418 => x"bb90528f",
   419 => x"51807270",
   420 => x"8405540c",
   421 => x"ff115170",
   422 => x"8025f238",
   423 => x"0288050d",
   424 => x"0402f005",
   425 => x"0d75518b",
   426 => x"e42d7082",
   427 => x"2cfc06bb",
   428 => x"90117210",
   429 => x"9e067108",
   430 => x"70722a70",
   431 => x"83068274",
   432 => x"2b700974",
   433 => x"06760c54",
   434 => x"51565753",
   435 => x"51538bde",
   436 => x"2d71bd9c",
   437 => x"0c029005",
   438 => x"0d0402fc",
   439 => x"050d7251",
   440 => x"80710c80",
   441 => x"0b84120c",
   442 => x"0284050d",
   443 => x"0402f005",
   444 => x"0d757008",
   445 => x"84120853",
   446 => x"5353ff54",
   447 => x"71712ea8",
   448 => x"388be42d",
   449 => x"84130870",
   450 => x"84291488",
   451 => x"11700870",
   452 => x"81ff0684",
   453 => x"18088111",
   454 => x"8706841a",
   455 => x"0c535155",
   456 => x"5151518b",
   457 => x"de2d7154",
   458 => x"73bd9c0c",
   459 => x"0290050d",
   460 => x"0402f805",
   461 => x"0d8be42d",
   462 => x"e008708b",
   463 => x"2a708106",
   464 => x"51525270",
   465 => x"802e9d38",
   466 => x"bdc40870",
   467 => x"8429bdcc",
   468 => x"057381ff",
   469 => x"06710c51",
   470 => x"51bdc408",
   471 => x"81118706",
   472 => x"bdc40c51",
   473 => x"800bbdec",
   474 => x"0c8bd72d",
   475 => x"8bde2d02",
   476 => x"88050d04",
   477 => x"02fc050d",
   478 => x"bdc4518d",
   479 => x"da2d8d84",
   480 => x"2d8eb151",
   481 => x"8bd32d02",
   482 => x"84050d04",
   483 => x"bdf008bd",
   484 => x"9c0c0402",
   485 => x"fc050d8f",
   486 => x"9d048bea",
   487 => x"2d80f651",
   488 => x"8da12dbd",
   489 => x"9c08f338",
   490 => x"80da518d",
   491 => x"a12dbd9c",
   492 => x"08e838bd",
   493 => x"9c08bbdc",
   494 => x"0cbd9c08",
   495 => x"5184f02d",
   496 => x"0284050d",
   497 => x"0402ec05",
   498 => x"0d765480",
   499 => x"52870b88",
   500 => x"1580f52d",
   501 => x"56537472",
   502 => x"248338a0",
   503 => x"53725182",
   504 => x"f92d8112",
   505 => x"8b1580f5",
   506 => x"2d545272",
   507 => x"7225de38",
   508 => x"0294050d",
   509 => x"0402f005",
   510 => x"0dbdf008",
   511 => x"5481f82d",
   512 => x"800bbdf4",
   513 => x"0c730880",
   514 => x"2e818038",
   515 => x"820bbdb0",
   516 => x"0cbdf408",
   517 => x"8f06bdac",
   518 => x"0c730852",
   519 => x"71832e96",
   520 => x"38718326",
   521 => x"89387181",
   522 => x"2eaf3890",
   523 => x"f6047185",
   524 => x"2e9f3890",
   525 => x"f6048814",
   526 => x"80f52d84",
   527 => x"1508b6f8",
   528 => x"53545285",
   529 => x"fe2d7184",
   530 => x"29137008",
   531 => x"525290fa",
   532 => x"0473518f",
   533 => x"c52d90f6",
   534 => x"04bbd808",
   535 => x"8815082c",
   536 => x"70810651",
   537 => x"5271802e",
   538 => x"8738b6fc",
   539 => x"5190f304",
   540 => x"b7805185",
   541 => x"fe2d8414",
   542 => x"085185fe",
   543 => x"2dbdf408",
   544 => x"8105bdf4",
   545 => x"0c8c1454",
   546 => x"90850402",
   547 => x"90050d04",
   548 => x"71bdf00c",
   549 => x"8ff52dbd",
   550 => x"f408ff05",
   551 => x"bdf80c04",
   552 => x"02e8050d",
   553 => x"bdf008bd",
   554 => x"fc085755",
   555 => x"87518da1",
   556 => x"2dbd9c08",
   557 => x"812a7081",
   558 => x"06515271",
   559 => x"802ea038",
   560 => x"91c6048b",
   561 => x"ea2d8751",
   562 => x"8da12dbd",
   563 => x"9c08f438",
   564 => x"bbdc0881",
   565 => x"3270bbdc",
   566 => x"0c705252",
   567 => x"84f02d80",
   568 => x"fe518da1",
   569 => x"2dbd9c08",
   570 => x"802ea638",
   571 => x"bbdc0880",
   572 => x"2e913880",
   573 => x"0bbbdc0c",
   574 => x"805184f0",
   575 => x"2d928304",
   576 => x"8bea2d80",
   577 => x"fe518da1",
   578 => x"2dbd9c08",
   579 => x"f33886e2",
   580 => x"2dbbdc08",
   581 => x"903881fd",
   582 => x"518da12d",
   583 => x"81fa518d",
   584 => x"a12d97d6",
   585 => x"0481f551",
   586 => x"8da12dbd",
   587 => x"9c08812a",
   588 => x"70810651",
   589 => x"5271802e",
   590 => x"af38bdf8",
   591 => x"08527180",
   592 => x"2e8938ff",
   593 => x"12bdf80c",
   594 => x"92e804bd",
   595 => x"f40810bd",
   596 => x"f4080570",
   597 => x"84291651",
   598 => x"52881208",
   599 => x"802e8938",
   600 => x"ff518812",
   601 => x"0852712d",
   602 => x"81f2518d",
   603 => x"a12dbd9c",
   604 => x"08812a70",
   605 => x"81065152",
   606 => x"71802eb1",
   607 => x"38bdf408",
   608 => x"ff11bdf8",
   609 => x"08565353",
   610 => x"73722589",
   611 => x"388114bd",
   612 => x"f80c93ad",
   613 => x"04721013",
   614 => x"70842916",
   615 => x"51528812",
   616 => x"08802e89",
   617 => x"38fe5188",
   618 => x"12085271",
   619 => x"2d81fd51",
   620 => x"8da12dbd",
   621 => x"9c08812a",
   622 => x"70810651",
   623 => x"5271802e",
   624 => x"ad38bdf8",
   625 => x"08802e89",
   626 => x"38800bbd",
   627 => x"f80c93ee",
   628 => x"04bdf408",
   629 => x"10bdf408",
   630 => x"05708429",
   631 => x"16515288",
   632 => x"1208802e",
   633 => x"8938fd51",
   634 => x"88120852",
   635 => x"712d81fa",
   636 => x"518da12d",
   637 => x"bd9c0881",
   638 => x"2a708106",
   639 => x"51527180",
   640 => x"2eae38bd",
   641 => x"f408ff11",
   642 => x"5452bdf8",
   643 => x"08732588",
   644 => x"3872bdf8",
   645 => x"0c94b004",
   646 => x"71101270",
   647 => x"84291651",
   648 => x"52881208",
   649 => x"802e8938",
   650 => x"fc518812",
   651 => x"0852712d",
   652 => x"bdf80870",
   653 => x"53547380",
   654 => x"2e8a388c",
   655 => x"15ff1555",
   656 => x"5594b604",
   657 => x"820bbdb0",
   658 => x"0c718f06",
   659 => x"bdac0c81",
   660 => x"eb518da1",
   661 => x"2dbd9c08",
   662 => x"812a7081",
   663 => x"06515271",
   664 => x"802ead38",
   665 => x"7408852e",
   666 => x"098106a4",
   667 => x"38881580",
   668 => x"f52dff05",
   669 => x"52718816",
   670 => x"81b72d71",
   671 => x"982b5271",
   672 => x"80258838",
   673 => x"800b8816",
   674 => x"81b72d74",
   675 => x"518fc52d",
   676 => x"81f4518d",
   677 => x"a12dbd9c",
   678 => x"08812a70",
   679 => x"81065152",
   680 => x"71802eb3",
   681 => x"38740885",
   682 => x"2e098106",
   683 => x"aa388815",
   684 => x"80f52d81",
   685 => x"05527188",
   686 => x"1681b72d",
   687 => x"7181ff06",
   688 => x"8b1680f5",
   689 => x"2d545272",
   690 => x"72278738",
   691 => x"72881681",
   692 => x"b72d7451",
   693 => x"8fc52d80",
   694 => x"da518da1",
   695 => x"2dbd9c08",
   696 => x"812a7081",
   697 => x"06515271",
   698 => x"802e81a6",
   699 => x"38bdf008",
   700 => x"bdf80855",
   701 => x"5373802e",
   702 => x"8a388c13",
   703 => x"ff155553",
   704 => x"95f50472",
   705 => x"08527182",
   706 => x"2ea63871",
   707 => x"82268938",
   708 => x"71812ea9",
   709 => x"38979204",
   710 => x"71832eb1",
   711 => x"3871842e",
   712 => x"09810680",
   713 => x"ed388813",
   714 => x"08519190",
   715 => x"2d979204",
   716 => x"bdf80851",
   717 => x"88130852",
   718 => x"712d9792",
   719 => x"04810b88",
   720 => x"14082bbb",
   721 => x"d80832bb",
   722 => x"d80c96e8",
   723 => x"04881380",
   724 => x"f52d8105",
   725 => x"8b1480f5",
   726 => x"2d535471",
   727 => x"74248338",
   728 => x"80547388",
   729 => x"1481b72d",
   730 => x"8ff52d97",
   731 => x"92047508",
   732 => x"802ea238",
   733 => x"7508518d",
   734 => x"a12dbd9c",
   735 => x"08810652",
   736 => x"71802e8b",
   737 => x"38bdf808",
   738 => x"51841608",
   739 => x"52712d88",
   740 => x"165675da",
   741 => x"38805480",
   742 => x"0bbdb00c",
   743 => x"738f06bd",
   744 => x"ac0ca052",
   745 => x"73bdf808",
   746 => x"2e098106",
   747 => x"9838bdf4",
   748 => x"08ff0574",
   749 => x"32700981",
   750 => x"05707207",
   751 => x"9f2a9171",
   752 => x"31515153",
   753 => x"53715182",
   754 => x"f92d8114",
   755 => x"548e7425",
   756 => x"c638bbdc",
   757 => x"085271bd",
   758 => x"9c0c0298",
   759 => x"050d0402",
   760 => x"f4050dd4",
   761 => x"5281ff72",
   762 => x"0c710853",
   763 => x"81ff720c",
   764 => x"72882b83",
   765 => x"fe800672",
   766 => x"087081ff",
   767 => x"06515253",
   768 => x"81ff720c",
   769 => x"72710788",
   770 => x"2b720870",
   771 => x"81ff0651",
   772 => x"525381ff",
   773 => x"720c7271",
   774 => x"07882b72",
   775 => x"087081ff",
   776 => x"067207bd",
   777 => x"9c0c5253",
   778 => x"028c050d",
   779 => x"0402f405",
   780 => x"0d747671",
   781 => x"81ff06d4",
   782 => x"0c5353be",
   783 => x"80088538",
   784 => x"71892b52",
   785 => x"71982ad4",
   786 => x"0c71902a",
   787 => x"7081ff06",
   788 => x"d40c5171",
   789 => x"882a7081",
   790 => x"ff06d40c",
   791 => x"517181ff",
   792 => x"06d40c72",
   793 => x"902a7081",
   794 => x"ff06d40c",
   795 => x"51d40870",
   796 => x"81ff0651",
   797 => x"5182b8bf",
   798 => x"527081ff",
   799 => x"2e098106",
   800 => x"943881ff",
   801 => x"0bd40cd4",
   802 => x"087081ff",
   803 => x"06ff1454",
   804 => x"515171e5",
   805 => x"3870bd9c",
   806 => x"0c028c05",
   807 => x"0d0402fc",
   808 => x"050d81c7",
   809 => x"5181ff0b",
   810 => x"d40cff11",
   811 => x"51708025",
   812 => x"f4380284",
   813 => x"050d0402",
   814 => x"f4050d81",
   815 => x"ff0bd40c",
   816 => x"93538052",
   817 => x"87fc80c1",
   818 => x"5198ad2d",
   819 => x"bd9c088b",
   820 => x"3881ff0b",
   821 => x"d40c8153",
   822 => x"99e40499",
   823 => x"9e2dff13",
   824 => x"5372df38",
   825 => x"72bd9c0c",
   826 => x"028c050d",
   827 => x"0402ec05",
   828 => x"0d810bbe",
   829 => x"800c8454",
   830 => x"d008708f",
   831 => x"2a708106",
   832 => x"51515372",
   833 => x"f33872d0",
   834 => x"0c999e2d",
   835 => x"b7845185",
   836 => x"fe2dd008",
   837 => x"708f2a70",
   838 => x"81065151",
   839 => x"5372f338",
   840 => x"810bd00c",
   841 => x"b1538052",
   842 => x"84d480c0",
   843 => x"5198ad2d",
   844 => x"bd9c0881",
   845 => x"2e933872",
   846 => x"822ebd38",
   847 => x"ff135372",
   848 => x"e538ff14",
   849 => x"5473ffb0",
   850 => x"38999e2d",
   851 => x"83aa5284",
   852 => x"9c80c851",
   853 => x"98ad2dbd",
   854 => x"9c08812e",
   855 => x"09810692",
   856 => x"3897df2d",
   857 => x"bd9c0883",
   858 => x"ffff0653",
   859 => x"7283aa2e",
   860 => x"9d3899b7",
   861 => x"2d9b8904",
   862 => x"b7905185",
   863 => x"fe2d8053",
   864 => x"9cd704b7",
   865 => x"a85185fe",
   866 => x"2d80549c",
   867 => x"a90481ff",
   868 => x"0bd40cb1",
   869 => x"54999e2d",
   870 => x"8fcf5380",
   871 => x"5287fc80",
   872 => x"f75198ad",
   873 => x"2dbd9c08",
   874 => x"55bd9c08",
   875 => x"812e0981",
   876 => x"069b3881",
   877 => x"ff0bd40c",
   878 => x"820a5284",
   879 => x"9c80e951",
   880 => x"98ad2dbd",
   881 => x"9c08802e",
   882 => x"8d38999e",
   883 => x"2dff1353",
   884 => x"72c9389c",
   885 => x"9c0481ff",
   886 => x"0bd40cbd",
   887 => x"9c085287",
   888 => x"fc80fa51",
   889 => x"98ad2dbd",
   890 => x"9c08b138",
   891 => x"81ff0bd4",
   892 => x"0cd40853",
   893 => x"81ff0bd4",
   894 => x"0c81ff0b",
   895 => x"d40c81ff",
   896 => x"0bd40c81",
   897 => x"ff0bd40c",
   898 => x"72862a70",
   899 => x"81067656",
   900 => x"51537295",
   901 => x"38bd9c08",
   902 => x"549ca904",
   903 => x"73822efe",
   904 => x"e238ff14",
   905 => x"5473feed",
   906 => x"3873be80",
   907 => x"0c738b38",
   908 => x"815287fc",
   909 => x"80d05198",
   910 => x"ad2d81ff",
   911 => x"0bd40cd0",
   912 => x"08708f2a",
   913 => x"70810651",
   914 => x"515372f3",
   915 => x"3872d00c",
   916 => x"81ff0bd4",
   917 => x"0c815372",
   918 => x"bd9c0c02",
   919 => x"94050d04",
   920 => x"02e8050d",
   921 => x"78558056",
   922 => x"81ff0bd4",
   923 => x"0cd00870",
   924 => x"8f2a7081",
   925 => x"06515153",
   926 => x"72f33882",
   927 => x"810bd00c",
   928 => x"81ff0bd4",
   929 => x"0c775287",
   930 => x"fc80d151",
   931 => x"98ad2d80",
   932 => x"dbc6df54",
   933 => x"bd9c0880",
   934 => x"2e8a38b7",
   935 => x"c85185fe",
   936 => x"2d9df704",
   937 => x"81ff0bd4",
   938 => x"0cd40870",
   939 => x"81ff0651",
   940 => x"537281fe",
   941 => x"2e098106",
   942 => x"9d3880ff",
   943 => x"5397df2d",
   944 => x"bd9c0875",
   945 => x"70840557",
   946 => x"0cff1353",
   947 => x"728025ed",
   948 => x"3881569d",
   949 => x"dc04ff14",
   950 => x"5473c938",
   951 => x"81ff0bd4",
   952 => x"0c81ff0b",
   953 => x"d40cd008",
   954 => x"708f2a70",
   955 => x"81065151",
   956 => x"5372f338",
   957 => x"72d00c75",
   958 => x"bd9c0c02",
   959 => x"98050d04",
   960 => x"02e8050d",
   961 => x"77797b58",
   962 => x"55558053",
   963 => x"727625a3",
   964 => x"38747081",
   965 => x"055680f5",
   966 => x"2d747081",
   967 => x"055680f5",
   968 => x"2d525271",
   969 => x"712e8638",
   970 => x"81519eb5",
   971 => x"04811353",
   972 => x"9e8c0480",
   973 => x"5170bd9c",
   974 => x"0c029805",
   975 => x"0d0402ec",
   976 => x"050d7655",
   977 => x"74802ebe",
   978 => x"389a1580",
   979 => x"e02d51ac",
   980 => x"822dbd9c",
   981 => x"08bd9c08",
   982 => x"80c4b40c",
   983 => x"bd9c0854",
   984 => x"5480c490",
   985 => x"08802e99",
   986 => x"38941580",
   987 => x"e02d51ac",
   988 => x"822dbd9c",
   989 => x"08902b83",
   990 => x"fff00a06",
   991 => x"70750751",
   992 => x"537280c4",
   993 => x"b40c80c4",
   994 => x"b4085372",
   995 => x"802e9d38",
   996 => x"80c48808",
   997 => x"fe147129",
   998 => x"80c49c08",
   999 => x"0580c4b8",
  1000 => x"0c70842b",
  1001 => x"80c4940c",
  1002 => x"549fda04",
  1003 => x"80c4a008",
  1004 => x"80c4b40c",
  1005 => x"80c4a408",
  1006 => x"80c4b80c",
  1007 => x"80c49008",
  1008 => x"802e8b38",
  1009 => x"80c48808",
  1010 => x"842b539f",
  1011 => x"d50480c4",
  1012 => x"a808842b",
  1013 => x"537280c4",
  1014 => x"940c0294",
  1015 => x"050d0402",
  1016 => x"d8050d80",
  1017 => x"0b80c490",
  1018 => x"0c845499",
  1019 => x"ed2dbd9c",
  1020 => x"08802e95",
  1021 => x"38be8452",
  1022 => x"80519ce0",
  1023 => x"2dbd9c08",
  1024 => x"802e8638",
  1025 => x"fe54a091",
  1026 => x"04ff1454",
  1027 => x"738024db",
  1028 => x"38738c38",
  1029 => x"b7d85185",
  1030 => x"fe2d7355",
  1031 => x"a5bb0480",
  1032 => x"56810b80",
  1033 => x"c4bc0c88",
  1034 => x"53b7ec52",
  1035 => x"beba519e",
  1036 => x"802dbd9c",
  1037 => x"08762e09",
  1038 => x"81068838",
  1039 => x"bd9c0880",
  1040 => x"c4bc0c88",
  1041 => x"53b7f852",
  1042 => x"bed6519e",
  1043 => x"802dbd9c",
  1044 => x"088838bd",
  1045 => x"9c0880c4",
  1046 => x"bc0c80c4",
  1047 => x"bc08802e",
  1048 => x"80fc3880",
  1049 => x"c1ca0b80",
  1050 => x"f52d80c1",
  1051 => x"cb0b80f5",
  1052 => x"2d71982b",
  1053 => x"71902b07",
  1054 => x"80c1cc0b",
  1055 => x"80f52d70",
  1056 => x"882b7207",
  1057 => x"80c1cd0b",
  1058 => x"80f52d71",
  1059 => x"0780c282",
  1060 => x"0b80f52d",
  1061 => x"80c2830b",
  1062 => x"80f52d71",
  1063 => x"882b0753",
  1064 => x"5f54525a",
  1065 => x"56575573",
  1066 => x"81abaa2e",
  1067 => x"0981068d",
  1068 => x"387551ab",
  1069 => x"d22dbd9c",
  1070 => x"0856a1ca",
  1071 => x"047382d4",
  1072 => x"d52e8738",
  1073 => x"b88451a2",
  1074 => x"8c04be84",
  1075 => x"5275519c",
  1076 => x"e02dbd9c",
  1077 => x"0855bd9c",
  1078 => x"08802e83",
  1079 => x"de388853",
  1080 => x"b7f852be",
  1081 => x"d6519e80",
  1082 => x"2dbd9c08",
  1083 => x"8a38810b",
  1084 => x"80c4900c",
  1085 => x"a2920488",
  1086 => x"53b7ec52",
  1087 => x"beba519e",
  1088 => x"802dbd9c",
  1089 => x"08802e8a",
  1090 => x"38b89851",
  1091 => x"85fe2da2",
  1092 => x"ee0480c2",
  1093 => x"820b80f5",
  1094 => x"2d547380",
  1095 => x"d52e0981",
  1096 => x"0680cb38",
  1097 => x"80c2830b",
  1098 => x"80f52d54",
  1099 => x"7381aa2e",
  1100 => x"098106ba",
  1101 => x"38800bbe",
  1102 => x"840b80f5",
  1103 => x"2d565474",
  1104 => x"81e92e83",
  1105 => x"38815474",
  1106 => x"81eb2e8c",
  1107 => x"38805573",
  1108 => x"752e0981",
  1109 => x"0682e438",
  1110 => x"be8f0b80",
  1111 => x"f52d5574",
  1112 => x"8d38be90",
  1113 => x"0b80f52d",
  1114 => x"5473822e",
  1115 => x"86388055",
  1116 => x"a5bb04be",
  1117 => x"910b80f5",
  1118 => x"2d7080c4",
  1119 => x"880cff05",
  1120 => x"80c48c0c",
  1121 => x"be920b80",
  1122 => x"f52dbe93",
  1123 => x"0b80f52d",
  1124 => x"58760577",
  1125 => x"82802905",
  1126 => x"7080c498",
  1127 => x"0cbe940b",
  1128 => x"80f52d70",
  1129 => x"80c4ac0c",
  1130 => x"80c49008",
  1131 => x"59575876",
  1132 => x"802e81ac",
  1133 => x"388853b7",
  1134 => x"f852bed6",
  1135 => x"519e802d",
  1136 => x"bd9c0881",
  1137 => x"f63880c4",
  1138 => x"88087084",
  1139 => x"2b80c494",
  1140 => x"0c7080c4",
  1141 => x"a80cbea9",
  1142 => x"0b80f52d",
  1143 => x"bea80b80",
  1144 => x"f52d7182",
  1145 => x"802905be",
  1146 => x"aa0b80f5",
  1147 => x"2d708480",
  1148 => x"802912be",
  1149 => x"ab0b80f5",
  1150 => x"2d708180",
  1151 => x"0a291270",
  1152 => x"80c4b00c",
  1153 => x"80c4ac08",
  1154 => x"712980c4",
  1155 => x"98080570",
  1156 => x"80c49c0c",
  1157 => x"beb10b80",
  1158 => x"f52dbeb0",
  1159 => x"0b80f52d",
  1160 => x"71828029",
  1161 => x"05beb20b",
  1162 => x"80f52d70",
  1163 => x"84808029",
  1164 => x"12beb30b",
  1165 => x"80f52d70",
  1166 => x"982b81f0",
  1167 => x"0a067205",
  1168 => x"7080c4a0",
  1169 => x"0cfe117e",
  1170 => x"29770580",
  1171 => x"c4a40c52",
  1172 => x"59524354",
  1173 => x"5e515259",
  1174 => x"525d5759",
  1175 => x"57a5b404",
  1176 => x"be960b80",
  1177 => x"f52dbe95",
  1178 => x"0b80f52d",
  1179 => x"71828029",
  1180 => x"057080c4",
  1181 => x"940c70a0",
  1182 => x"2983ff05",
  1183 => x"70892a70",
  1184 => x"80c4a80c",
  1185 => x"be9b0b80",
  1186 => x"f52dbe9a",
  1187 => x"0b80f52d",
  1188 => x"71828029",
  1189 => x"057080c4",
  1190 => x"b00c7b71",
  1191 => x"291e7080",
  1192 => x"c4a40c7d",
  1193 => x"80c4a00c",
  1194 => x"730580c4",
  1195 => x"9c0c555e",
  1196 => x"51515555",
  1197 => x"80519ebe",
  1198 => x"2d815574",
  1199 => x"bd9c0c02",
  1200 => x"a8050d04",
  1201 => x"02ec050d",
  1202 => x"7670872c",
  1203 => x"7180ff06",
  1204 => x"55565480",
  1205 => x"c490088a",
  1206 => x"3873882c",
  1207 => x"7481ff06",
  1208 => x"5455be84",
  1209 => x"5280c498",
  1210 => x"0815519c",
  1211 => x"e02dbd9c",
  1212 => x"0854bd9c",
  1213 => x"08802eb4",
  1214 => x"3880c490",
  1215 => x"08802e98",
  1216 => x"38728429",
  1217 => x"be840570",
  1218 => x"085253ab",
  1219 => x"d22dbd9c",
  1220 => x"08f00a06",
  1221 => x"53a6aa04",
  1222 => x"7210be84",
  1223 => x"057080e0",
  1224 => x"2d5253ac",
  1225 => x"822dbd9c",
  1226 => x"08537254",
  1227 => x"73bd9c0c",
  1228 => x"0294050d",
  1229 => x"0402e005",
  1230 => x"0d797084",
  1231 => x"2c80c4b8",
  1232 => x"0805718f",
  1233 => x"06525553",
  1234 => x"728938be",
  1235 => x"84527351",
  1236 => x"9ce02d72",
  1237 => x"a029be84",
  1238 => x"05548074",
  1239 => x"80f52d56",
  1240 => x"5374732e",
  1241 => x"83388153",
  1242 => x"7481e52e",
  1243 => x"81f13881",
  1244 => x"70740654",
  1245 => x"5872802e",
  1246 => x"81e5388b",
  1247 => x"1480f52d",
  1248 => x"70832a79",
  1249 => x"06585676",
  1250 => x"9938bbe0",
  1251 => x"08537289",
  1252 => x"387280c2",
  1253 => x"840b81b7",
  1254 => x"2d76bbe0",
  1255 => x"0c7353a8",
  1256 => x"e104758f",
  1257 => x"2e098106",
  1258 => x"81b53874",
  1259 => x"9f068d29",
  1260 => x"80c1f711",
  1261 => x"51538114",
  1262 => x"80f52d73",
  1263 => x"70810555",
  1264 => x"81b72d83",
  1265 => x"1480f52d",
  1266 => x"73708105",
  1267 => x"5581b72d",
  1268 => x"851480f5",
  1269 => x"2d737081",
  1270 => x"055581b7",
  1271 => x"2d871480",
  1272 => x"f52d7370",
  1273 => x"81055581",
  1274 => x"b72d8914",
  1275 => x"80f52d73",
  1276 => x"70810555",
  1277 => x"81b72d8e",
  1278 => x"1480f52d",
  1279 => x"73708105",
  1280 => x"5581b72d",
  1281 => x"901480f5",
  1282 => x"2d737081",
  1283 => x"055581b7",
  1284 => x"2d921480",
  1285 => x"f52d7370",
  1286 => x"81055581",
  1287 => x"b72d9414",
  1288 => x"80f52d73",
  1289 => x"70810555",
  1290 => x"81b72d96",
  1291 => x"1480f52d",
  1292 => x"73708105",
  1293 => x"5581b72d",
  1294 => x"981480f5",
  1295 => x"2d737081",
  1296 => x"055581b7",
  1297 => x"2d9c1480",
  1298 => x"f52d7370",
  1299 => x"81055581",
  1300 => x"b72d9e14",
  1301 => x"80f52d73",
  1302 => x"81b72d77",
  1303 => x"bbe00c80",
  1304 => x"5372bd9c",
  1305 => x"0c02a005",
  1306 => x"0d0402cc",
  1307 => x"050d7e60",
  1308 => x"5e5a800b",
  1309 => x"80c4b408",
  1310 => x"80c4b808",
  1311 => x"595c5680",
  1312 => x"5880c494",
  1313 => x"08782e81",
  1314 => x"b038778f",
  1315 => x"06a01757",
  1316 => x"54738f38",
  1317 => x"be845276",
  1318 => x"51811757",
  1319 => x"9ce02dbe",
  1320 => x"84568076",
  1321 => x"80f52d56",
  1322 => x"5474742e",
  1323 => x"83388154",
  1324 => x"7481e52e",
  1325 => x"80f73881",
  1326 => x"70750655",
  1327 => x"5c73802e",
  1328 => x"80eb388b",
  1329 => x"1680f52d",
  1330 => x"98065978",
  1331 => x"80df388b",
  1332 => x"537c5275",
  1333 => x"519e802d",
  1334 => x"bd9c0880",
  1335 => x"d0389c16",
  1336 => x"0851abd2",
  1337 => x"2dbd9c08",
  1338 => x"841b0c9a",
  1339 => x"1680e02d",
  1340 => x"51ac822d",
  1341 => x"bd9c08bd",
  1342 => x"9c08881c",
  1343 => x"0cbd9c08",
  1344 => x"555580c4",
  1345 => x"9008802e",
  1346 => x"98389416",
  1347 => x"80e02d51",
  1348 => x"ac822dbd",
  1349 => x"9c08902b",
  1350 => x"83fff00a",
  1351 => x"06701651",
  1352 => x"5473881b",
  1353 => x"0c787a0c",
  1354 => x"7b54aaf2",
  1355 => x"04811858",
  1356 => x"80c49408",
  1357 => x"7826fed2",
  1358 => x"3880c490",
  1359 => x"08802eb0",
  1360 => x"387a51a5",
  1361 => x"c42dbd9c",
  1362 => x"08bd9c08",
  1363 => x"80ffffff",
  1364 => x"f806555b",
  1365 => x"7380ffff",
  1366 => x"fff82e94",
  1367 => x"38bd9c08",
  1368 => x"fe0580c4",
  1369 => x"88082980",
  1370 => x"c49c0805",
  1371 => x"57a8ff04",
  1372 => x"805473bd",
  1373 => x"9c0c02b4",
  1374 => x"050d0402",
  1375 => x"f4050d74",
  1376 => x"70088105",
  1377 => x"710c7008",
  1378 => x"80c48c08",
  1379 => x"06535371",
  1380 => x"8e388813",
  1381 => x"0851a5c4",
  1382 => x"2dbd9c08",
  1383 => x"88140c81",
  1384 => x"0bbd9c0c",
  1385 => x"028c050d",
  1386 => x"0402f005",
  1387 => x"0d758811",
  1388 => x"08fe0580",
  1389 => x"c4880829",
  1390 => x"80c49c08",
  1391 => x"11720880",
  1392 => x"c48c0806",
  1393 => x"05795553",
  1394 => x"54549ce0",
  1395 => x"2d029005",
  1396 => x"0d0402f4",
  1397 => x"050d7470",
  1398 => x"882a83fe",
  1399 => x"80067072",
  1400 => x"982a0772",
  1401 => x"882b87fc",
  1402 => x"80800673",
  1403 => x"982b81f0",
  1404 => x"0a067173",
  1405 => x"0707bd9c",
  1406 => x"0c565153",
  1407 => x"51028c05",
  1408 => x"0d0402f8",
  1409 => x"050d028e",
  1410 => x"0580f52d",
  1411 => x"74882b07",
  1412 => x"7083ffff",
  1413 => x"06bd9c0c",
  1414 => x"51028805",
  1415 => x"0d0402f4",
  1416 => x"050d7476",
  1417 => x"78535452",
  1418 => x"80712597",
  1419 => x"38727081",
  1420 => x"055480f5",
  1421 => x"2d727081",
  1422 => x"055481b7",
  1423 => x"2dff1151",
  1424 => x"70eb3880",
  1425 => x"7281b72d",
  1426 => x"028c050d",
  1427 => x"0402e805",
  1428 => x"0d775680",
  1429 => x"70565473",
  1430 => x"7624b338",
  1431 => x"80c49408",
  1432 => x"742eab38",
  1433 => x"7351a6b5",
  1434 => x"2dbd9c08",
  1435 => x"bd9c0809",
  1436 => x"810570bd",
  1437 => x"9c08079f",
  1438 => x"2a770581",
  1439 => x"17575753",
  1440 => x"53747624",
  1441 => x"893880c4",
  1442 => x"94087426",
  1443 => x"d73872bd",
  1444 => x"9c0c0298",
  1445 => x"050d0402",
  1446 => x"f0050dbd",
  1447 => x"98081651",
  1448 => x"accd2dbd",
  1449 => x"9c08802e",
  1450 => x"9e388b53",
  1451 => x"bd9c0852",
  1452 => x"80c28451",
  1453 => x"ac9e2d80",
  1454 => x"c4c00854",
  1455 => x"73802e87",
  1456 => x"3880c284",
  1457 => x"51732d02",
  1458 => x"90050d04",
  1459 => x"02dc050d",
  1460 => x"80705a55",
  1461 => x"74bd9808",
  1462 => x"25b13880",
  1463 => x"c4940875",
  1464 => x"2ea93878",
  1465 => x"51a6b52d",
  1466 => x"bd9c0809",
  1467 => x"810570bd",
  1468 => x"9c08079f",
  1469 => x"2a760581",
  1470 => x"1b5b5654",
  1471 => x"74bd9808",
  1472 => x"25893880",
  1473 => x"c4940879",
  1474 => x"26d93880",
  1475 => x"557880c4",
  1476 => x"94082781",
  1477 => x"d4387851",
  1478 => x"a6b52dbd",
  1479 => x"9c08802e",
  1480 => x"81a838bd",
  1481 => x"9c088b05",
  1482 => x"80f52d70",
  1483 => x"842a7081",
  1484 => x"06771078",
  1485 => x"842b80c2",
  1486 => x"840b80f5",
  1487 => x"2d5c5c53",
  1488 => x"51555673",
  1489 => x"802e80c9",
  1490 => x"38741682",
  1491 => x"2bb08d0b",
  1492 => x"bbec120c",
  1493 => x"54777531",
  1494 => x"1080c4c4",
  1495 => x"11555690",
  1496 => x"74708105",
  1497 => x"5681b72d",
  1498 => x"a07481b7",
  1499 => x"2d7681ff",
  1500 => x"06811658",
  1501 => x"5473802e",
  1502 => x"8a389c53",
  1503 => x"80c28452",
  1504 => x"af89048b",
  1505 => x"53bd9c08",
  1506 => x"5280c4c6",
  1507 => x"1651afc2",
  1508 => x"04741682",
  1509 => x"2bad970b",
  1510 => x"bbec120c",
  1511 => x"547681ff",
  1512 => x"06811658",
  1513 => x"5473802e",
  1514 => x"8a389c53",
  1515 => x"80c28452",
  1516 => x"afb9048b",
  1517 => x"53bd9c08",
  1518 => x"52777531",
  1519 => x"1080c4c4",
  1520 => x"05517655",
  1521 => x"ac9e2daf",
  1522 => x"de047490",
  1523 => x"29753170",
  1524 => x"1080c4c4",
  1525 => x"055154bd",
  1526 => x"9c087481",
  1527 => x"b72d8119",
  1528 => x"59748b24",
  1529 => x"a338ae8d",
  1530 => x"04749029",
  1531 => x"75317010",
  1532 => x"80c4c405",
  1533 => x"8c773157",
  1534 => x"51548074",
  1535 => x"81b72d9e",
  1536 => x"14ff1656",
  1537 => x"5474f338",
  1538 => x"02a4050d",
  1539 => x"0402fc05",
  1540 => x"0dbd9808",
  1541 => x"1351accd",
  1542 => x"2dbd9c08",
  1543 => x"802e8838",
  1544 => x"bd9c0851",
  1545 => x"9ebe2d80",
  1546 => x"0bbd980c",
  1547 => x"adcc2d8f",
  1548 => x"f52d0284",
  1549 => x"050d0402",
  1550 => x"fc050d72",
  1551 => x"5170fd2e",
  1552 => x"ad3870fd",
  1553 => x"248a3870",
  1554 => x"fc2e80c4",
  1555 => x"38b19804",
  1556 => x"70fe2eb1",
  1557 => x"3870ff2e",
  1558 => x"098106bc",
  1559 => x"38bd9808",
  1560 => x"5170802e",
  1561 => x"b338ff11",
  1562 => x"bd980cb1",
  1563 => x"9804bd98",
  1564 => x"08f00570",
  1565 => x"bd980c51",
  1566 => x"7080259c",
  1567 => x"38800bbd",
  1568 => x"980cb198",
  1569 => x"04bd9808",
  1570 => x"8105bd98",
  1571 => x"0cb19804",
  1572 => x"bd980890",
  1573 => x"05bd980c",
  1574 => x"adcc2d8f",
  1575 => x"f52d0284",
  1576 => x"050d0402",
  1577 => x"fc050d80",
  1578 => x"0bbd980c",
  1579 => x"adcc2d8f",
  1580 => x"8c2dbd9c",
  1581 => x"08bd880c",
  1582 => x"bbe45191",
  1583 => x"902d0284",
  1584 => x"050d0471",
  1585 => x"80c4c00c",
  1586 => x"04000000",
  1587 => x"00ffffff",
  1588 => x"ff00ffff",
  1589 => x"ffff00ff",
  1590 => x"ffffff00",
  1591 => x"52657365",
  1592 => x"74000000",
  1593 => x"43617267",
  1594 => x"61722044",
  1595 => x"6973636f",
  1596 => x"2f43696e",
  1597 => x"74612010",
  1598 => x"00000000",
  1599 => x"45786974",
  1600 => x"00000000",
  1601 => x"46444320",
  1602 => x"4f726967",
  1603 => x"696e616c",
  1604 => x"00000000",
  1605 => x"46444320",
  1606 => x"46617374",
  1607 => x"00000000",
  1608 => x"4d756c74",
  1609 => x"69666163",
  1610 => x"65203220",
  1611 => x"456e6162",
  1612 => x"6c656400",
  1613 => x"4d756c74",
  1614 => x"69666163",
  1615 => x"65203220",
  1616 => x"48696464",
  1617 => x"656e0000",
  1618 => x"4d756c74",
  1619 => x"69666163",
  1620 => x"65203220",
  1621 => x"44697361",
  1622 => x"626c6564",
  1623 => x"00000000",
  1624 => x"4d6f7573",
  1625 => x"65204469",
  1626 => x"7361626c",
  1627 => x"65640000",
  1628 => x"4d6f7573",
  1629 => x"6520456e",
  1630 => x"61626c65",
  1631 => x"64000000",
  1632 => x"506c6179",
  1633 => x"63697479",
  1634 => x"20446973",
  1635 => x"61626c65",
  1636 => x"64000000",
  1637 => x"506c6179",
  1638 => x"63697479",
  1639 => x"20456e61",
  1640 => x"626c6564",
  1641 => x"00000000",
  1642 => x"52696768",
  1643 => x"74205368",
  1644 => x"69667420",
  1645 => x"61732042",
  1646 => x"61636b73",
  1647 => x"6c617368",
  1648 => x"00000000",
  1649 => x"52696768",
  1650 => x"74205368",
  1651 => x"69667420",
  1652 => x"61732053",
  1653 => x"68696674",
  1654 => x"00000000",
  1655 => x"536f756e",
  1656 => x"64206f75",
  1657 => x"74707574",
  1658 => x"20537465",
  1659 => x"72656f00",
  1660 => x"536f756e",
  1661 => x"64206f75",
  1662 => x"74707574",
  1663 => x"204d6f6e",
  1664 => x"6f000000",
  1665 => x"54617065",
  1666 => x"20736f75",
  1667 => x"6e642044",
  1668 => x"69736162",
  1669 => x"6c656400",
  1670 => x"54617065",
  1671 => x"20736f75",
  1672 => x"6e642045",
  1673 => x"6e61626c",
  1674 => x"65640000",
  1675 => x"43505520",
  1676 => x"74696d69",
  1677 => x"6e677320",
  1678 => x"4f726967",
  1679 => x"696e616c",
  1680 => x"00000000",
  1681 => x"43505520",
  1682 => x"74696d69",
  1683 => x"6e677320",
  1684 => x"46617374",
  1685 => x"00000000",
  1686 => x"53696e63",
  1687 => x"20736967",
  1688 => x"6e616c73",
  1689 => x"204f7269",
  1690 => x"67696e61",
  1691 => x"6c000000",
  1692 => x"53696e63",
  1693 => x"20736967",
  1694 => x"6e616c73",
  1695 => x"2046696c",
  1696 => x"74657265",
  1697 => x"64000000",
  1698 => x"43525443",
  1699 => x"20547970",
  1700 => x"65203100",
  1701 => x"43525443",
  1702 => x"20547970",
  1703 => x"65203200",
  1704 => x"44697370",
  1705 => x"6c617920",
  1706 => x"436f6c6f",
  1707 => x"72284741",
  1708 => x"29000000",
  1709 => x"44697370",
  1710 => x"6c617920",
  1711 => x"436f6c6f",
  1712 => x"72202841",
  1713 => x"53494329",
  1714 => x"00000000",
  1715 => x"44697370",
  1716 => x"6c617920",
  1717 => x"47726565",
  1718 => x"6e000000",
  1719 => x"44697370",
  1720 => x"6c617920",
  1721 => x"416d6265",
  1722 => x"72000000",
  1723 => x"44697370",
  1724 => x"6c617920",
  1725 => x"4379616e",
  1726 => x"00000000",
  1727 => x"44697370",
  1728 => x"6c617920",
  1729 => x"57686974",
  1730 => x"65000000",
  1731 => x"5363616e",
  1732 => x"6c696e65",
  1733 => x"73204e6f",
  1734 => x"6e650000",
  1735 => x"5363616e",
  1736 => x"6c696e65",
  1737 => x"73204352",
  1738 => x"54203235",
  1739 => x"25000000",
  1740 => x"5363616e",
  1741 => x"6c696e65",
  1742 => x"73204352",
  1743 => x"54203530",
  1744 => x"25000000",
  1745 => x"5363616e",
  1746 => x"6c696e65",
  1747 => x"73204352",
  1748 => x"54203735",
  1749 => x"25000000",
  1750 => x"43617267",
  1751 => x"61204661",
  1752 => x"6c6c6964",
  1753 => x"61000000",
  1754 => x"4f4b0000",
  1755 => x"414d5354",
  1756 => x"52414420",
  1757 => x"44415400",
  1758 => x"16200000",
  1759 => x"14200000",
  1760 => x"15200000",
  1761 => x"53442069",
  1762 => x"6e69742e",
  1763 => x"2e2e0a00",
  1764 => x"53442063",
  1765 => x"61726420",
  1766 => x"72657365",
  1767 => x"74206661",
  1768 => x"696c6564",
  1769 => x"210a0000",
  1770 => x"53444843",
  1771 => x"20657272",
  1772 => x"6f72210a",
  1773 => x"00000000",
  1774 => x"57726974",
  1775 => x"65206661",
  1776 => x"696c6564",
  1777 => x"0a000000",
  1778 => x"52656164",
  1779 => x"20666169",
  1780 => x"6c65640a",
  1781 => x"00000000",
  1782 => x"43617264",
  1783 => x"20696e69",
  1784 => x"74206661",
  1785 => x"696c6564",
  1786 => x"0a000000",
  1787 => x"46415431",
  1788 => x"36202020",
  1789 => x"00000000",
  1790 => x"46415433",
  1791 => x"32202020",
  1792 => x"00000000",
  1793 => x"4e6f2070",
  1794 => x"61727469",
  1795 => x"74696f6e",
  1796 => x"20736967",
  1797 => x"0a000000",
  1798 => x"42616420",
  1799 => x"70617274",
  1800 => x"0a000000",
  1801 => x"4261636b",
  1802 => x"00000000",
  1803 => x"00000002",
  1804 => x"00000002",
  1805 => x"000018dc",
  1806 => x"0000034e",
  1807 => x"00000003",
  1808 => x"00001d5c",
  1809 => x"00000004",
  1810 => x"00000003",
  1811 => x"00001d44",
  1812 => x"00000006",
  1813 => x"00000003",
  1814 => x"00001d3c",
  1815 => x"00000002",
  1816 => x"00000003",
  1817 => x"00001d34",
  1818 => x"00000002",
  1819 => x"00000003",
  1820 => x"00001d2c",
  1821 => x"00000002",
  1822 => x"00000003",
  1823 => x"00001d24",
  1824 => x"00000002",
  1825 => x"00000003",
  1826 => x"00001d1c",
  1827 => x"00000002",
  1828 => x"00000003",
  1829 => x"00001d14",
  1830 => x"00000002",
  1831 => x"00000003",
  1832 => x"00001d0c",
  1833 => x"00000002",
  1834 => x"00000003",
  1835 => x"00001d04",
  1836 => x"00000002",
  1837 => x"00000003",
  1838 => x"00001cf8",
  1839 => x"00000003",
  1840 => x"00000003",
  1841 => x"00001cf0",
  1842 => x"00000002",
  1843 => x"00000002",
  1844 => x"000018e4",
  1845 => x"000018a3",
  1846 => x"00000002",
  1847 => x"000018fc",
  1848 => x"00000793",
  1849 => x"00000000",
  1850 => x"00000000",
  1851 => x"00000000",
  1852 => x"00001904",
  1853 => x"00001914",
  1854 => x"00001920",
  1855 => x"00001934",
  1856 => x"00001948",
  1857 => x"00001960",
  1858 => x"00001970",
  1859 => x"00001980",
  1860 => x"00001994",
  1861 => x"000019a8",
  1862 => x"000019c4",
  1863 => x"000019dc",
  1864 => x"000019f0",
  1865 => x"00001a04",
  1866 => x"00001a18",
  1867 => x"00001a2c",
  1868 => x"00001a44",
  1869 => x"00001a58",
  1870 => x"00001a70",
  1871 => x"00001a88",
  1872 => x"00001a94",
  1873 => x"00001aa0",
  1874 => x"00001ab4",
  1875 => x"00001acc",
  1876 => x"00001adc",
  1877 => x"00001aec",
  1878 => x"00001afc",
  1879 => x"00001b0c",
  1880 => x"00001b1c",
  1881 => x"00001b30",
  1882 => x"00001b44",
  1883 => x"00000004",
  1884 => x"00001b58",
  1885 => x"00001d6c",
  1886 => x"00000004",
  1887 => x"00001b68",
  1888 => x"00001c30",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"00000000",
  1894 => x"00000000",
  1895 => x"00000000",
  1896 => x"00000000",
  1897 => x"00000000",
  1898 => x"00000000",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000002",
  1914 => x"00002244",
  1915 => x"00001697",
  1916 => x"00000002",
  1917 => x"00002262",
  1918 => x"00001697",
  1919 => x"00000002",
  1920 => x"00002280",
  1921 => x"00001697",
  1922 => x"00000002",
  1923 => x"0000229e",
  1924 => x"00001697",
  1925 => x"00000002",
  1926 => x"000022bc",
  1927 => x"00001697",
  1928 => x"00000002",
  1929 => x"000022da",
  1930 => x"00001697",
  1931 => x"00000002",
  1932 => x"000022f8",
  1933 => x"00001697",
  1934 => x"00000002",
  1935 => x"00002316",
  1936 => x"00001697",
  1937 => x"00000002",
  1938 => x"00002334",
  1939 => x"00001697",
  1940 => x"00000002",
  1941 => x"00002352",
  1942 => x"00001697",
  1943 => x"00000002",
  1944 => x"00002370",
  1945 => x"00001697",
  1946 => x"00000002",
  1947 => x"0000238e",
  1948 => x"00001697",
  1949 => x"00000002",
  1950 => x"000023ac",
  1951 => x"00001697",
  1952 => x"00000004",
  1953 => x"00001c24",
  1954 => x"00000000",
  1955 => x"00000000",
  1956 => x"00000000",
  1957 => x"00001837",
  1958 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

